--------------------------------------------------------------
-- Project          : VHDL description of ARC processor (chapter 5)
--                    "Computer Architecture and Organisation" (ISBN 978-0-471-73388-1) by Murdocca and Heuring
-- 
-- File             : main_memory_arch.vhd
--
-- Related File(s)  : conversion_utilites.vhd
--
-- Author           : E. Molenkamp, University of Twente, the Netherlands
-- Email            : e.molenkamp@utwente.nl
-- 
-- Project          : Computer Organization
-- Creation Date    : 27 June 2008
-- 
-- Contents         : Architecure of main memory.
--                    Memory is filled with bin filegenerated by the ARCtools  
--                    (default for program is  "program.bin"; see entity main_memory) .
--
-- Change Log 
--   Author         : E.Molenkamp
--   Email          : e.molenkamp@utwente.nl
--   Date           : 16 October 2008 
--   Changes        : Function fill_memory is changed in an IMPURE function
--
ARCHITECTURE bhv OF main_memory IS

  TYPE mem_tp IS ARRAY (0 TO max_address/4-1) OF string(1 TO 8);
    
  IMPURE FUNCTION fill_memory (program : string) RETURN mem_tp IS
    VARIABLE mem : mem_tp := (OTHERS=>(OTHERS=>'-'));
    FILE prg : text OPEN read_mode IS program;
    VARIABLE inp_line : line;
    VARIABLE str : string(1 TO 8);
    VARIABLE addr : natural;
	VARIABLE char : character;
  BEGIN
    READLINE(prg, inp_line); -- the first line in the BIN file generated by the ARCTOOLS is to be ignored
    WHILE NOT endfile(prg) LOOP
      READLINE(prg,inp_line);
      READ(inp_line, str); -- address is read;
      addr := hex2dec(str);
	  ASSERT (addr MOD 4)=0 REPORT "address not multiple of 4" SEVERITY error;
      READ(inp_line,char); -- read TAB
      READ(inp_line, str); -- 
      mem(addr/4):=str;
    END LOOP;
	RETURN mem;
  END fill_memory;
  
  SIGNAL mem : mem_tp := fill_memory(program);   

BEGIN
  
  
  ACK <= '1'; -- it is assmued that the memory can deliver the data within one cycle
  
  PROCESS (clk)
  BEGIN
    IF falling_edge(clk) THEN
      IF Wr_M='1' THEN
        ASSERT address(1 DOWNTO 0)="00" REPORT "write to main memory: not aligned address (should be multiple of 4)" SEVERITY warning;	  
        mem(to_integer(unsigned(address(31 downto 2)))) <= stdv2hexv(DataIn);
      END IF;  
    END IF;
  END PROCESS;

  -- The address bus is connected with the A bus. Hence not all data on the A bus is
  -- used as an address. It could be out of the implemented address range.
  Dout <= hexv2stdv(mem(to_integer(unsigned(address(31 downto 2))))) WHEN Rd_M='1' ELSE
          (OTHERS=>'-'); -- word addressing

  ASSERT (Rd_M='1' AND address(1 DOWNTO 0)="00") OR (Rd_M/='1')
    REPORT "read from main memory: not aligned address (should be multiple of 4)" SEVERITY warning;		  
		  
END bhv;

